// tests that use and test private functions
module time